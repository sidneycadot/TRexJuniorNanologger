
package constants is

    constant NUM_INPUTS : positive := 8;

    constant SAMPLE_BITS_PER_CLOCK : positive := 8;

    constant FIFO_WIDTH : positive := 117;
    constant FIFO_DEPTH : positive := 8192;

end package constants;
